// ===============================
// RISCV_Single_Cycle.v (Đã sửa)
// ===============================

module RISCV_Single_Cycle (
    input clk,
    input rst_n,
    output [31:0] PC_out_top,
    output [31:0] Instruction_out_top,
    output [31:0] x[0:31],
    output [31:0] dmem[0:255]
);

    // Wires
    wire [31:0] pc_out, pc_in, inst, imm, read_data1, read_data2, alu_result, mem_read_data, write_data;
    wire [31:0] alu_operand2, pc_plus_4, branch_target, jalr_target;
    wire reg_write, mem_read, mem_write, mem_to_reg, alu_src, branch, jump, zero;
    wire [3:0] alu_op;
    wire [1:0] pc_src;
    wire pc_write;

    // PC logic
    assign pc_write = 1'b1;
    assign pc_plus_4 = pc_out + 4;
    assign branch_target = pc_out + imm;
    assign jalr_target = read_data1 + imm;
    assign pc_in = (pc_src == 2'b00) ? pc_plus_4 :
                   (pc_src == 2'b01) ? branch_target :
                   (pc_src == 2'b10) ? jalr_target : pc_plus_4;

    PC pc_inst (
        .clk(clk),
        .rst_n(rst_n),
        .pc_in(pc_in),
        .pc_write(pc_write),
        .pc_out(pc_out)
    );

    // IMEM
    IMEM IMEM_inst (
        .addr(pc_out),
        .inst(inst)
    );

    // Control Unit
    ControlUnit ctrl_inst (
        .opcode(inst[6:0]),
        .funct3(inst[14:12]),
        .funct7(inst[31:25]),
        .reg_write(reg_write),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .mem_to_reg(mem_to_reg),
        .alu_op(alu_op),
        .alu_src(alu_src),
        .branch(branch),
        .jump(jump),
        .pc_src(pc_src)
    );

    // Register File
    RegisterFile Reg_inst (
        .clk(clk),
        .rst_n(rst_n),
        .rs1(inst[19:15]),
        .rs2(inst[24:20]),
        .rd(inst[11:7]),
        .write_data(write_data),
        .reg_write(reg_write),
        .read_data1(read_data1),
        .read_data2(read_data2)
    );

    // Immediate Generator
    ImmGen imm_gen_inst (
        .inst(inst),
        .imm(imm)
    );

    // ALU
    assign alu_operand2 = alu_src ? imm : read_data2;
    ALU alu_inst (
        .operand1(read_data1),
        .operand2(alu_operand2),
        .alu_op(alu_op),
        .result(alu_result),
        .zero(zero)
    );

    // Data Memory
    DMEM DMEM_inst (
        .clk(clk),
        .addr(alu_result),
        .write_data(read_data2),
        .mem_write(mem_write),
        .mem_read(mem_read),
        .read_data(mem_read_data)
    );

    // Write-back
    assign write_data = mem_to_reg ? mem_read_data : 
                        (jump ? pc_plus_4 : alu_result);

    // Outputs for testbench
    assign PC_out_top = pc_out;
    assign Instruction_out_top = inst;

    genvar i;
    generate
        for (i = 0; i < 32; i = i + 1) begin
            assign x[i] = Reg_inst.registers[i];
        end
        for (i = 0; i < 256; i = i + 1) begin
            assign dmem[i] = DMEM_inst.memory[i];
        end
    endgenerate
endmodule
